module fourBitAdder_tb;
    reg A[3:0],B[3:0],Cin;
    wire S[3:0],Cout;
    initial begin
        $dum
        A = 4'b0001;
    end

endmodule