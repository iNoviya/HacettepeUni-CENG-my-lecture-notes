`timescale 1 ns/10 ps
module full_adder_tb;


endmodule